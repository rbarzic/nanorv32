module GNDPAD (/*AUTOARG*/);

   

   /*AUTOINPUT*/
   /*AUTOOUTPUT*/

   /*AUTOREG*/
   /*AUTOWIRE*/

endmodule // GNDPAD
/*
 Local Variables:
 verilog-library-directories:(
 "."
 )
 End:
 */
