module rfiniocell (/*AUTOARG*/
   // Outputs
   rfin,
   // Inouts
   PAD
   );

   inout wire  PAD;

   output wire rfin;
   
   
   /*AUTOINPUT*/
   /*AUTOOUTPUT*/

   /*AUTOREG*/
   /*AUTOWIRE*/

   assign rfin = PAD;
   
endmodule // rfiniocell
/*
 Local Variables:
 verilog-library-directories:(
 "."
 )
 End:
 */
