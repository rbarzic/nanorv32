module CORNER;

   

   /*AUTOREG*/
   /*AUTOWIRE*/

endmodule // CORNER
/*
 Local Variables:
 verilog-library-directories:(
 "."
 )
 End:
 */
