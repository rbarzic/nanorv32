module ESDPAD (/*AUTOARG*/);

   

   /*AUTOINPUT*/
   /*AUTOOUTPUT*/

   /*AUTOREG*/
   /*AUTOWIRE*/

endmodule // ESDPAD
/*
 Local Variables:
 verilog-library-directories:(
 "."
 )
 End:
 */
