module PWRPAD (/*AUTOARG*/);

   

   /*AUTOINPUT*/
   /*AUTOOUTPUT*/

   /*AUTOREG*/
   /*AUTOWIRE*/

endmodule // PWRPAD
/*
 Local Variables:
 verilog-library-directories:(
 "."
 )
 End:
 */
