VERSION 5.6 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;

MACRO bytewrite_ram_32bits
    CLASS BLOCK ;
    FOREIGN bytewrite_ram_32bits 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 150.0 BY 300.0 ;
    SYMMETRY x y r90 ;

    PIN dvcc
        DIRECTION  INOUT ;
	USE POWER ;
        PORT
        LAYER MET1 ;
        RECT  46.8 295.2 51.6 300.0 ;
        END
    END dvcc

    PIN dgnd
        DIRECTION  INOUT ;
	USE GROUND ;
        PORT
        LAYER MET1 ;
        RECT  98.4 295.2 103.2 300.0 ;
        END
    END dgnd

    PIN dout[0]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 8.76 150.0 9.0 ;
        END
    END dout[0]

    PIN dout[1]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 17.76 150.0 18.0 ;
        END
    END dout[1]

    PIN dout[2]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 26.76 150.0 27.0 ;
        END
    END dout[2]

    PIN dout[3]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 35.76 150.0 36.0 ;
        END
    END dout[3]

    PIN dout[4]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 44.76 150.0 45.0 ;
        END
    END dout[4]

    PIN dout[5]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 53.76 150.0 54.0 ;
        END
    END dout[5]

    PIN dout[6]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 62.76 150.0 63.0 ;
        END
    END dout[6]

    PIN dout[7]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 71.76 150.0 72.0 ;
        END
    END dout[7]

    PIN dout[8]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 80.76 150.0 81.0 ;
        END
    END dout[8]

    PIN dout[9]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 89.76 150.0 90.0 ;
        END
    END dout[9]

    PIN dout[10]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 98.76 150.0 99.0 ;
        END
    END dout[10]

    PIN dout[11]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 107.76 150.0 108.0 ;
        END
    END dout[11]

    PIN dout[12]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 116.76 150.0 117.0 ;
        END
    END dout[12]

    PIN dout[13]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 125.76 150.0 126.0 ;
        END
    END dout[13]

    PIN dout[14]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 134.76 150.0 135.0 ;
        END
    END dout[14]

    PIN dout[15]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 143.76 150.0 144.0 ;
        END
    END dout[15]

    PIN dout[16]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 152.76 150.0 153.0 ;
        END
    END dout[16]

    PIN dout[17]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 161.76 150.0 162.0 ;
        END
    END dout[17]

    PIN dout[18]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 170.76 150.0 171.0 ;
        END
    END dout[18]

    PIN dout[19]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 179.76 150.0 180.0 ;
        END
    END dout[19]

    PIN dout[20]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 188.76 150.0 189.0 ;
        END
    END dout[20]

    PIN dout[21]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 197.76 150.0 198.0 ;
        END
    END dout[21]

    PIN dout[22]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 206.76 150.0 207.0 ;
        END
    END dout[22]

    PIN dout[23]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 215.76 150.0 216.0 ;
        END
    END dout[23]

    PIN dout[24]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 224.76 150.0 225.0 ;
        END
    END dout[24]

    PIN dout[25]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 233.76 150.0 234.0 ;
        END
    END dout[25]

    PIN dout[26]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 242.76 150.0 243.0 ;
        END
    END dout[26]

    PIN dout[27]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 251.76 150.0 252.0 ;
        END
    END dout[27]

    PIN dout[28]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 260.76 150.0 261.0 ;
        END
    END dout[28]

    PIN dout[29]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 269.76 150.0 270.0 ;
        END
    END dout[29]

    PIN dout[30]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 278.76 150.0 279.0 ;
        END
    END dout[30]

    PIN dout[31]
        DIRECTION  OUTPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  149.76 287.76 150.0 288.0 ;
        END
    END dout[31]

    PIN clk
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 5.76 0.24 6.0 ;
        END
    END clk

    PIN we[0]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 11.76 0.24 12.0 ;
        END
    END we[0]

    PIN we[1]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 17.76 0.24 18.0 ;
        END
    END we[1]

    PIN we[2]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 23.76 0.24 24.0 ;
        END
    END we[2]

    PIN we[3]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 29.76 0.24 30.0 ;
        END
    END we[3]

    PIN din[0]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 35.76 0.24 36.0 ;
        END
    END din[0]

    PIN din[1]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 41.76 0.24 42.0 ;
        END
    END din[1]

    PIN din[2]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 47.76 0.24 48.0 ;
        END
    END din[2]

    PIN din[3]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 53.76 0.24 54.0 ;
        END
    END din[3]

    PIN din[4]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 59.76 0.24 60.0 ;
        END
    END din[4]

    PIN din[5]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 65.76 0.24 66.0 ;
        END
    END din[5]

    PIN din[6]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 71.76 0.24 72.0 ;
        END
    END din[6]

    PIN din[7]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 77.76 0.24 78.0 ;
        END
    END din[7]

    PIN din[8]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 83.76 0.24 84.0 ;
        END
    END din[8]

    PIN din[9]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 89.76 0.24 90.0 ;
        END
    END din[9]

    PIN din[10]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 95.76 0.24 96.0 ;
        END
    END din[10]

    PIN din[11]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 101.76 0.24 102.0 ;
        END
    END din[11]

    PIN din[12]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 107.76 0.24 108.0 ;
        END
    END din[12]

    PIN din[13]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 113.76 0.24 114.0 ;
        END
    END din[13]

    PIN din[14]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 119.76 0.24 120.0 ;
        END
    END din[14]

    PIN din[15]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 125.76 0.24 126.0 ;
        END
    END din[15]

    PIN din[16]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 131.76 0.24 132.0 ;
        END
    END din[16]

    PIN din[17]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 137.76 0.24 138.0 ;
        END
    END din[17]

    PIN din[18]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 143.76 0.24 144.0 ;
        END
    END din[18]

    PIN din[19]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 149.76 0.24 150.0 ;
        END
    END din[19]

    PIN din[20]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 155.76 0.24 156.0 ;
        END
    END din[20]

    PIN din[21]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 161.76 0.24 162.0 ;
        END
    END din[21]

    PIN din[22]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 167.76 0.24 168.0 ;
        END
    END din[22]

    PIN din[23]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 173.76 0.24 174.0 ;
        END
    END din[23]

    PIN din[24]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 179.76 0.24 180.0 ;
        END
    END din[24]

    PIN din[25]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 185.76 0.24 186.0 ;
        END
    END din[25]

    PIN din[26]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 191.76 0.24 192.0 ;
        END
    END din[26]

    PIN din[27]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 197.76 0.24 198.0 ;
        END
    END din[27]

    PIN din[28]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 203.76 0.24 204.0 ;
        END
    END din[28]

    PIN din[29]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 209.76 0.24 210.0 ;
        END
    END din[29]

    PIN din[30]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 215.76 0.24 216.0 ;
        END
    END din[30]

    PIN din[31]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 221.76 0.24 222.0 ;
        END
    END din[31]

    PIN addr[0]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 227.76 0.24 228.0 ;
        END
    END addr[0]

    PIN addr[1]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 233.76 0.24 234.0 ;
        END
    END addr[1]

    PIN addr[2]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 239.76 0.24 240.0 ;
        END
    END addr[2]

    PIN addr[3]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 245.76 0.24 246.0 ;
        END
    END addr[3]

    PIN addr[4]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 251.76 0.24 252.0 ;
        END
    END addr[4]

    PIN addr[5]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 257.76 0.24 258.0 ;
        END
    END addr[5]

    PIN addr[6]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 263.76 0.24 264.0 ;
        END
    END addr[6]

    PIN addr[7]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 269.76 0.24 270.0 ;
        END
    END addr[7]

    PIN addr[8]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 275.76 0.24 276.0 ;
        END
    END addr[8]

    PIN addr[9]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 281.76 0.24 282.0 ;
        END
    END addr[9]

    PIN addr[10]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 287.76 0.24 288.0 ;
        END
    END addr[10]

    PIN addr[11]
        DIRECTION  INPUT ;
	
        PORT
        LAYER MET1 ;
        RECT  0 293.76 0.24 294.0 ;
        END
    END addr[11]

END bytewrite_ram_32bits

END LIBRARY
