module anaiocell (/*AUTOARG*/
   // Outputs
   ao18in,
   // Inouts
   PAD
   );

   inout wire  PAD;

   output wire ao18in;
   

   /*AUTOINPUT*/
   /*AUTOOUTPUT*/

   /*AUTOREG*/
   /*AUTOWIRE*/

   assign ao18in = PAD;
endmodule // anaiocell
/*
 Local Variables:
 verilog-library-directories:(
 "."
 )
 End:
 */
