/*
  *  PicoRV32 -- A Small RISC-V (RV32I) Processor Core
  *
  *  Copyright (C) 2015  Clifford Wolf <clifford@clifford.at>
  *
  *  Permission to use, copy, modify, and/or distribute this software for any
  *  purpose with or without fee is hereby granted, provided that the above
  *  copyright notice and this permission notice appear in all copies.
  *
  *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
  *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
  *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
  *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
  *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
  *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
  *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
  *
  */

`timescale 1 ns / 1 ps
  // `default_nettype none
  // `define DEBUG

`ifdef DEBUG
 `define debug(debug_command) debug_command
`else
 `define debug(debug_command)
`endif

`ifdef FORMAL
 `define FORMAL_KEEP (* keep *)
`else
 `define FORMAL_KEEP
`endif

  /***************************************************************
   * picorv32
   ***************************************************************/

  module picorv32 #(
                    parameter [ 0:0] ENABLE_COUNTERS = 1,
	            parameter [ 0:0] ENABLE_REGS_16_31 = 1,
	            parameter [ 0:0] ENABLE_REGS_DUALPORT = 1,
	            parameter [ 0:0] LATCHED_MEM_RDATA = 0,
	            parameter [ 0:0] TWO_STAGE_SHIFT = 1,
	            parameter [ 0:0] TWO_CYCLE_COMPARE = 0,
	            parameter [ 0:0] TWO_CYCLE_ALU = 0,
	            parameter [ 0:0] CATCH_MISALIGN = 1,
	            parameter [ 0:0] CATCH_ILLINSN = 1,
	            parameter [ 0:0] ENABLE_PCPI = 0,
	            parameter [ 0:0] ENABLE_MUL = 0,
	            parameter [ 0:0] ENABLE_IRQ = 0,
	            parameter [ 0:0] ENABLE_IRQ_QREGS = 1,
	            parameter [ 0:0] ENABLE_IRQ_TIMER = 1,
	            parameter [31:0] MASKED_IRQ = 32'h 0000_0000,
	            parameter [31:0] LATCHED_IRQ = 32'h ffff_ffff,
	            parameter [31:0] PROGADDR_RESET = 32'h 0000_0000,
	            parameter [31:0] PROGADDR_IRQ = 32'h 0000_0010
                    ) (
	               input             clk, resetn,
	               output reg        trap,

	               output reg        mem_valid,
	               output reg        mem_instr,
	               input             mem_ready,

	               output reg [31:0] mem_addr,
	               output reg [31:0] mem_wdata,
	               output reg [ 3:0] mem_wstrb,
	               input [31:0]      mem_rdata,

	               // Look-Ahead Interface
	               output            mem_la_read,
	               output            mem_la_write,
	               output [31:0]     mem_la_addr,
	               output reg [31:0] mem_la_wdata,
	               output reg [ 3:0] mem_la_wstrb,

	               // Pico Co-Processor Interface (PCPI)
	               output reg        pcpi_valid,
	               output reg [31:0] pcpi_insn,
	               output [31:0]     pcpi_rs1,
	               output [31:0]     pcpi_rs2,
	               input             pcpi_wr,
	               input [31:0]      pcpi_rd,
	               input             pcpi_wait,
	               input             pcpi_ready,

	               // IRQ Interface
	               input [31:0]      irq,
	               output reg [31:0] eoi
                       );
   localparam integer                    irq_timer = 0;
   localparam integer                    irq_sbreak = 1;
   localparam integer                    irq_buserror = 2;

   localparam integer                    irqregs_offset = ENABLE_REGS_16_31 ? 32 : 16;
   localparam integer                    regfile_size = (ENABLE_REGS_16_31 ? 32 : 16) + 4*ENABLE_IRQ*ENABLE_IRQ_QREGS;
   localparam integer                    regindex_bits = (ENABLE_REGS_16_31 ? 5 : 4) + ENABLE_IRQ*ENABLE_IRQ_QREGS;

   localparam WITH_PCPI = ENABLE_PCPI || ENABLE_MUL;

   reg [63:0]                            count_cycle, count_instr;
   reg [31:0]                            reg_pc, reg_next_pc, reg_op1, reg_op2, reg_out;
   reg [31:0]                            cpuregs [0:regfile_size-1];
   reg [4:0]                             reg_sh;

   assign pcpi_rs1 = reg_op1;
   assign pcpi_rs2 = reg_op2;

   wire [31:0]                           next_pc;

   reg                                   irq_active;
   reg [31:0]                            irq_mask;
   reg [31:0]                            irq_pending;
   reg [31:0]                            timer;


   // Internal PCPI Cores

   wire                                  pcpi_mul_wr;
   wire [31:0]                           pcpi_mul_rd;
   wire                                  pcpi_mul_wait;
   wire                                  pcpi_mul_ready;

   reg                                   pcpi_int_wr;
   reg [31:0]                            pcpi_int_rd;
   reg                                   pcpi_int_wait;
   reg                                   pcpi_int_ready;


   wire [31:0]                           x0,x1,x2,x3,x4,x5,x6,x7;
   wire [31:0]                           a0,a1,a2,a3,a4,a5,a6,a7;
   assign x0 = cpuregs[0];
   assign x1 = cpuregs[1];
   assign x2 = cpuregs[2];
   assign x3 = cpuregs[3];
   assign x4 = cpuregs[4];
   assign x5 = cpuregs[5];
   assign x6 = cpuregs[6];
   assign x7 = cpuregs[7];


   assign a0 = cpuregs[18];
   assign a1 = cpuregs[19];
   assign a2 = cpuregs[20];
   assign a3 = cpuregs[21];
   assign a4 = cpuregs[22];
   assign a5 = cpuregs[23];
   assign a6 = cpuregs[24];
   assign a7 = cpuregs[25];



   generate if (ENABLE_MUL) begin
      picorv32_pcpi_mul pcpi_mul (
			          .clk       (clk            ),
			          .resetn    (resetn         ),
			          .pcpi_valid(pcpi_valid     ),
			          .pcpi_insn (pcpi_insn      ),
			          .pcpi_rs1  (pcpi_rs1       ),
			          .pcpi_rs2  (pcpi_rs2       ),
			          .pcpi_wr   (pcpi_mul_wr    ),
			          .pcpi_rd   (pcpi_mul_rd    ),
			          .pcpi_wait (pcpi_mul_wait  ),
			          .pcpi_ready(pcpi_mul_ready )
		                  );
   end else begin
      assign pcpi_mul_wr = 0;
      assign pcpi_mul_rd = 1'bx;
      assign pcpi_mul_wait = 0;
      assign pcpi_mul_ready = 0;
   end endgenerate

   always @* begin
      pcpi_int_wr = 0;
      pcpi_int_rd = 1'bx;
      pcpi_int_wait  = |{ENABLE_PCPI && pcpi_wait,  ENABLE_MUL && pcpi_mul_wait};
      pcpi_int_ready = |{ENABLE_PCPI && pcpi_ready, ENABLE_MUL && pcpi_mul_ready};

      (* parallel_case *)
      case (1'b1)
	ENABLE_PCPI && pcpi_ready: begin
	   pcpi_int_wr = pcpi_wr;
	   pcpi_int_rd = pcpi_rd;
	end
	ENABLE_MUL && pcpi_mul_ready: begin
	   pcpi_int_wr = pcpi_mul_wr;
	   pcpi_int_rd = pcpi_mul_rd;
	end
      endcase
   end


   // Memory Interface

   reg [1:0] mem_state;
   reg [1:0] mem_wordsize;
   reg [31:0] mem_rdata_word;
   reg [31:0] mem_rdata_q;
   reg        mem_do_prefetch;
   reg        mem_do_rinst;
   reg        mem_do_rdata;
   reg        mem_do_wdata;

   wire       mem_busy = |{mem_do_prefetch, mem_do_rinst, mem_do_rdata, mem_do_wdata};
   wire       mem_done = resetn && ((mem_ready && |mem_state && (mem_do_rinst || mem_do_rdata || mem_do_wdata)) || (&mem_state && mem_do_rinst));

   assign mem_la_write = resetn && !mem_state && mem_do_wdata;
   assign mem_la_read = resetn && !mem_state && (mem_do_rinst || mem_do_prefetch || mem_do_rdata);
   assign mem_la_addr = (mem_do_prefetch || mem_do_rinst) ? next_pc : {reg_op1[31:2], 2'b00};

   wire [31:0] mem_rdata_latched;
   assign mem_rdata_latched = ((mem_valid && mem_ready) || LATCHED_MEM_RDATA) ? mem_rdata : mem_rdata_q;

   always @* begin
      (* full_case *)
      case (mem_wordsize)
	0: begin
	   mem_la_wdata = reg_op2;
	   mem_la_wstrb = 4'b1111;
	   mem_rdata_word = mem_rdata;
	end
	1: begin
	   mem_la_wdata = {2{reg_op2[15:0]}};
	   mem_la_wstrb = reg_op1[1] ? 4'b1100 : 4'b0011;
	   case (reg_op1[1])
	     1'b0: mem_rdata_word = mem_rdata[15: 0];
	     1'b1: mem_rdata_word = mem_rdata[31:16];
	   endcase
	end
	2: begin
	   mem_la_wdata = {4{reg_op2[7:0]}};
	   mem_la_wstrb = 4'b0001 << reg_op1[1:0];
	   case (reg_op1[1:0])
	     2'b00: mem_rdata_word = mem_rdata[ 7: 0];
	     2'b01: mem_rdata_word = mem_rdata[15: 8];
	     2'b10: mem_rdata_word = mem_rdata[23:16];
	     2'b11: mem_rdata_word = mem_rdata[31:24];
	   endcase
	end
      endcase
   end

   always @(posedge clk) begin
      if (mem_valid && mem_ready)
	mem_rdata_q <= mem_rdata_latched;
   end

   always @(posedge clk) begin
      if (!resetn) begin
	 mem_state <= 0;
	 mem_valid <= 0;
      end else case (mem_state)
		 0: begin
		    mem_addr <= mem_la_addr;
		    mem_wdata <= mem_la_wdata;
		    mem_wstrb <= mem_la_wstrb;
		    if (mem_do_prefetch || mem_do_rinst || mem_do_rdata) begin
		       mem_valid <= 1;
		       mem_instr <= mem_do_prefetch || mem_do_rinst;
		       mem_wstrb <= 0;
		       mem_state <= 1;
		    end
		    if (mem_do_wdata) begin
		       mem_valid <= 1;
		       mem_instr <= 0;
		       mem_state <= 2;
		    end
		 end
		 1: begin
		    if (mem_ready) begin
		       mem_valid <= 0;
		       mem_state <= mem_do_rinst || mem_do_rdata ? 0 : 3;
		    end
		 end
		 2: begin
		    if (mem_ready) begin
		       mem_valid <= 0;
		       mem_state <= 0;
		    end
		 end
		 3: begin
		    if (mem_do_rinst) begin
		       mem_state <= 0;
		    end
		 end
	       endcase
   end


   // Instruction Decoder

   reg instr_lui, instr_auipc, instr_jal, instr_jalr;
   reg instr_beq, instr_bne, instr_blt, instr_bge, instr_bltu, instr_bgeu;
   reg instr_lb, instr_lh, instr_lw, instr_lbu, instr_lhu, instr_sb, instr_sh, instr_sw;
   reg instr_addi, instr_slti, instr_sltiu, instr_xori, instr_ori, instr_andi, instr_slli, instr_srli, instr_srai;
   reg instr_add, instr_sub, instr_sll, instr_slt, instr_sltu, instr_xor, instr_srl, instr_sra, instr_or, instr_and;
   reg instr_rdcycle, instr_rdcycleh, instr_rdinstr, instr_rdinstrh;
   reg instr_getq, instr_setq, instr_retirq, instr_maskirq, instr_waitirq, instr_timer;
   wire instr_trap;

   reg [regindex_bits-1:0] decoded_rd, decoded_rs1, decoded_rs2;
   reg [31:0]              decoded_imm, decoded_imm_uj;
   reg                     decoder_trigger;
   reg                     decoder_trigger_q;
   reg                     decoder_pseudo_trigger;

   reg                     is_lui_auipc_jal;
   reg                     is_lb_lh_lw_lbu_lhu;
   reg                     is_slli_srli_srai;
   reg                     is_jalr_addi_slti_sltiu_xori_ori_andi;
   reg                     is_sb_sh_sw;
   reg                     is_sll_srl_sra;
   reg                     is_lui_auipc_jal_jalr_addi_add_sub;
   reg                     is_slti_blt_slt;
   reg                     is_sltiu_bltu_sltu;
   reg                     is_beq_bne_blt_bge_bltu_bgeu;
   reg                     is_lbu_lhu_lw;
   reg                     is_alu_reg_imm;
   reg                     is_alu_reg_reg;
   reg                     is_compare;

   assign instr_trap = (CATCH_ILLINSN || ENABLE_PCPI) && !{instr_lui, instr_auipc, instr_jal, instr_jalr,
			                                   instr_beq, instr_bne, instr_blt, instr_bge, instr_bltu, instr_bgeu,
			                                   instr_lb, instr_lh, instr_lw, instr_lbu, instr_lhu, instr_sb, instr_sh, instr_sw,
			                                   instr_addi, instr_slti, instr_sltiu, instr_xori, instr_ori, instr_andi, instr_slli, instr_srli, instr_srai,
			                                   instr_add, instr_sub, instr_sll, instr_slt, instr_sltu, instr_xor, instr_srl, instr_sra, instr_or, instr_and,
			                                   instr_rdcycle, instr_rdcycleh, instr_rdinstr, instr_rdinstrh,
			                                   instr_getq, instr_setq, instr_retirq, instr_maskirq, instr_waitirq, instr_timer};

   wire                    is_rdcycle_rdcycleh_rdinstr_rdinstrh;
   assign is_rdcycle_rdcycleh_rdinstr_rdinstrh = |{instr_rdcycle, instr_rdcycleh, instr_rdinstr, instr_rdinstrh};

   reg [63:0]              new_ascii_instr;
   `FORMAL_KEEP reg [63:0] ascii_instr;

   always @(posedge clk) begin
      new_ascii_instr = "";
      if (instr_lui)      new_ascii_instr = "lui";
      if (instr_auipc)    new_ascii_instr = "auipc";
      if (instr_jal)      new_ascii_instr = "jal";
      if (instr_jalr)     new_ascii_instr = "jalr";

      if (instr_beq)      new_ascii_instr = "beq";
      if (instr_bne)      new_ascii_instr = "bne";
      if (instr_blt)      new_ascii_instr = "blt";
      if (instr_bge)      new_ascii_instr = "bge";
      if (instr_bltu)     new_ascii_instr = "bltu";
      if (instr_bgeu)     new_ascii_instr = "bgeu";

      if (instr_lb)       new_ascii_instr = "lb";
      if (instr_lh)       new_ascii_instr = "lh";
      if (instr_lw)       new_ascii_instr = "lw";
      if (instr_lbu)      new_ascii_instr = "lbu";
      if (instr_lhu)      new_ascii_instr = "lhu";
      if (instr_sb)       new_ascii_instr = "sb";
      if (instr_sh)       new_ascii_instr = "sh";
      if (instr_sw)       new_ascii_instr = "sw";

      if (instr_addi)     new_ascii_instr = "addi";
      if (instr_slti)     new_ascii_instr = "slti";
      if (instr_sltiu)    new_ascii_instr = "sltiu";
      if (instr_xori)     new_ascii_instr = "xori";
      if (instr_ori)      new_ascii_instr = "ori";
      if (instr_andi)     new_ascii_instr = "andi";
      if (instr_slli)     new_ascii_instr = "slli";
      if (instr_srli)     new_ascii_instr = "srli";
      if (instr_srai)     new_ascii_instr = "srai";

      if (instr_add)      new_ascii_instr = "add";
      if (instr_sub)      new_ascii_instr = "sub";
      if (instr_sll)      new_ascii_instr = "sll";
      if (instr_slt)      new_ascii_instr = "slt";
      if (instr_sltu)     new_ascii_instr = "sltu";
      if (instr_xor)      new_ascii_instr = "xor";
      if (instr_srl)      new_ascii_instr = "srl";
      if (instr_sra)      new_ascii_instr = "sra";
      if (instr_or)       new_ascii_instr = "or";
      if (instr_and)      new_ascii_instr = "and";

      if (instr_rdcycle)  new_ascii_instr = "rdcycle";
      if (instr_rdcycleh) new_ascii_instr = "rdcycleh";
      if (instr_rdinstr)  new_ascii_instr = "rdinstr";
      if (instr_rdinstrh) new_ascii_instr = "rdinstrh";

      if (instr_getq)     new_ascii_instr = "getq";
      if (instr_setq)     new_ascii_instr = "setq";
      if (instr_retirq)   new_ascii_instr = "retirq";
      if (instr_maskirq)  new_ascii_instr = "maskirq";
      if (instr_waitirq)  new_ascii_instr = "waitirq";
      if (instr_timer)    new_ascii_instr = "timer";

      if (decoder_trigger_q)
	ascii_instr <= new_ascii_instr;
   end

   always @(posedge clk) begin
      is_lui_auipc_jal <= |{instr_lui, instr_auipc, instr_jal};
      is_lui_auipc_jal_jalr_addi_add_sub <= |{instr_lui, instr_auipc, instr_jal, instr_jalr, instr_addi, instr_add, instr_sub};
      is_slti_blt_slt <= |{instr_slti, instr_blt, instr_slt};
      is_sltiu_bltu_sltu <= |{instr_sltiu, instr_bltu, instr_sltu};
      is_lbu_lhu_lw <= |{instr_lbu, instr_lhu, instr_lw};
      is_compare <= |{is_beq_bne_blt_bge_bltu_bgeu, instr_slti, instr_slt, instr_sltiu, instr_sltu};

      if (mem_do_rinst && mem_done) begin
	 instr_lui     <= mem_rdata_latched[6:0] == 7'b0110111;
	 instr_auipc   <= mem_rdata_latched[6:0] == 7'b0010111;
	 instr_jal     <= mem_rdata_latched[6:0] == 7'b1101111;
	 instr_jalr    <= mem_rdata_latched[6:0] == 7'b1100111;
	 instr_retirq  <= mem_rdata_latched[6:0] == 7'b0001011 && mem_rdata_latched[31:25] == 7'b0000010 && ENABLE_IRQ;
	 instr_waitirq <= mem_rdata_latched[6:0] == 7'b0001011 && mem_rdata_latched[31:25] == 7'b0000100 && ENABLE_IRQ;

	 is_beq_bne_blt_bge_bltu_bgeu <= mem_rdata_latched[6:0] == 7'b1100011;
	 is_lb_lh_lw_lbu_lhu          <= mem_rdata_latched[6:0] == 7'b0000011;
	 is_sb_sh_sw                  <= mem_rdata_latched[6:0] == 7'b0100011;
	 is_alu_reg_imm               <= mem_rdata_latched[6:0] == 7'b0010011;
	 is_alu_reg_reg               <= mem_rdata_latched[6:0] == 7'b0110011;

	 { decoded_imm_uj[31:20], decoded_imm_uj[10:1], decoded_imm_uj[11], decoded_imm_uj[19:12], decoded_imm_uj[0] } <= $signed({mem_rdata_latched[31:12], 1'b0});

	 decoded_rd <= mem_rdata_latched[11:7];
	 decoded_rs1 <= mem_rdata_latched[19:15];
	 decoded_rs2 <= mem_rdata_latched[24:20];

	 if (mem_rdata_latched[6:0] == 7'b0001011 && mem_rdata_latched[31:25] == 7'b0000000 && ENABLE_IRQ && ENABLE_IRQ_QREGS)
	   decoded_rs1[regindex_bits-1] <= 1; // instr_getq

	 if (mem_rdata_latched[6:0] == 7'b0001011 && mem_rdata_latched[31:25] == 7'b0000010 && ENABLE_IRQ)
	   decoded_rs1 <= ENABLE_IRQ_QREGS ? irqregs_offset : 3; // instr_retirq
      end

      if (decoder_trigger && !decoder_pseudo_trigger) begin
	 pcpi_insn <= WITH_PCPI ? mem_rdata_q : 'bx;

	 instr_beq   <= is_beq_bne_blt_bge_bltu_bgeu && mem_rdata_q[14:12] == 3'b000;
	 instr_bne   <= is_beq_bne_blt_bge_bltu_bgeu && mem_rdata_q[14:12] == 3'b001;
	 instr_blt   <= is_beq_bne_blt_bge_bltu_bgeu && mem_rdata_q[14:12] == 3'b100;
	 instr_bge   <= is_beq_bne_blt_bge_bltu_bgeu && mem_rdata_q[14:12] == 3'b101;
	 instr_bltu  <= is_beq_bne_blt_bge_bltu_bgeu && mem_rdata_q[14:12] == 3'b110;
	 instr_bgeu  <= is_beq_bne_blt_bge_bltu_bgeu && mem_rdata_q[14:12] == 3'b111;

	 instr_lb    <= is_lb_lh_lw_lbu_lhu && mem_rdata_q[14:12] == 3'b000;
	 instr_lh    <= is_lb_lh_lw_lbu_lhu && mem_rdata_q[14:12] == 3'b001;
	 instr_lw    <= is_lb_lh_lw_lbu_lhu && mem_rdata_q[14:12] == 3'b010;
	 instr_lbu   <= is_lb_lh_lw_lbu_lhu && mem_rdata_q[14:12] == 3'b100;
	 instr_lhu   <= is_lb_lh_lw_lbu_lhu && mem_rdata_q[14:12] == 3'b101;

	 instr_sb    <= is_sb_sh_sw && mem_rdata_q[14:12] == 3'b000;
	 instr_sh    <= is_sb_sh_sw && mem_rdata_q[14:12] == 3'b001;
	 instr_sw    <= is_sb_sh_sw && mem_rdata_q[14:12] == 3'b010;

	 instr_addi  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b000;
	 instr_slti  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b010;
	 instr_sltiu <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b011;
	 instr_xori  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b100;
	 instr_ori   <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b110;
	 instr_andi  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b111;

	 instr_slli  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b001 && mem_rdata_q[31:25] == 7'b0000000;
	 instr_srli  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0000000;
	 instr_srai  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0100000;

	 instr_add   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b000 && mem_rdata_q[31:25] == 7'b0000000;
	 instr_sub   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b000 && mem_rdata_q[31:25] == 7'b0100000;
	 instr_sll   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b001 && mem_rdata_q[31:25] == 7'b0000000;
	 instr_slt   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b010 && mem_rdata_q[31:25] == 7'b0000000;
	 instr_sltu  <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b011 && mem_rdata_q[31:25] == 7'b0000000;
	 instr_xor   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b100 && mem_rdata_q[31:25] == 7'b0000000;
	 instr_srl   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0000000;
	 instr_sra   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0100000;
	 instr_or    <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b110 && mem_rdata_q[31:25] == 7'b0000000;
	 instr_and   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b111 && mem_rdata_q[31:25] == 7'b0000000;

	 instr_rdcycle  <= ((mem_rdata_q[6:0] == 7'b1110011 && mem_rdata_q[31:12] == 'b11000000000000000010) ||
			    (mem_rdata_q[6:0] == 7'b1110011 && mem_rdata_q[31:12] == 'b11000000000100000010)) && ENABLE_COUNTERS;
	 instr_rdcycleh <= ((mem_rdata_q[6:0] == 7'b1110011 && mem_rdata_q[31:12] == 'b11001000000000000010) ||
			    (mem_rdata_q[6:0] == 7'b1110011 && mem_rdata_q[31:12] == 'b11001000000100000010)) && ENABLE_COUNTERS;
	 instr_rdinstr  <=  (mem_rdata_q[6:0] == 7'b1110011 && mem_rdata_q[31:12] == 'b11000000001000000010) && ENABLE_COUNTERS;
	 instr_rdinstrh <=  (mem_rdata_q[6:0] == 7'b1110011 && mem_rdata_q[31:12] == 'b11001000001000000010) && ENABLE_COUNTERS;

	 instr_getq    <= mem_rdata_q[6:0] == 7'b0001011 && mem_rdata_q[31:25] == 7'b0000000 && ENABLE_IRQ && ENABLE_IRQ_QREGS;
	 instr_setq    <= mem_rdata_q[6:0] == 7'b0001011 && mem_rdata_q[31:25] == 7'b0000001 && ENABLE_IRQ && ENABLE_IRQ_QREGS;
	 instr_maskirq <= mem_rdata_q[6:0] == 7'b0001011 && mem_rdata_q[31:25] == 7'b0000011 && ENABLE_IRQ;
	 instr_timer   <= mem_rdata_q[6:0] == 7'b0001011 && mem_rdata_q[31:25] == 7'b0000101 && ENABLE_IRQ && ENABLE_IRQ_TIMER;

	 is_slli_srli_srai <= is_alu_reg_imm && |{
				                  mem_rdata_q[14:12] == 3'b001 && mem_rdata_q[31:25] == 7'b0000000,
				                  mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0000000,
				                  mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0100000
			                          };

	 is_jalr_addi_slti_sltiu_xori_ori_andi <= instr_jalr || is_alu_reg_imm && |{
				                                                    mem_rdata_q[14:12] == 3'b000,
				                                                    mem_rdata_q[14:12] == 3'b010,
				                                                    mem_rdata_q[14:12] == 3'b011,
				                                                    mem_rdata_q[14:12] == 3'b100,
				                                                    mem_rdata_q[14:12] == 3'b110,
				                                                    mem_rdata_q[14:12] == 3'b111
			                                                            };

	 is_sll_srl_sra <= is_alu_reg_reg && |{
				               mem_rdata_q[14:12] == 3'b001 && mem_rdata_q[31:25] == 7'b0000000,
				               mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0000000,
				               mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0100000
			                       };

	 (* parallel_case *)
	 case (1'b1)
	   instr_jal:
	     decoded_imm <= decoded_imm_uj;
	   |{instr_lui, instr_auipc}:
			    decoded_imm <= mem_rdata_q[31:12] << 12;
	   |{instr_jalr, is_lb_lh_lw_lbu_lhu, is_alu_reg_imm}:
			    decoded_imm <= $signed(mem_rdata_q[31:20]);
	   is_beq_bne_blt_bge_bltu_bgeu:
	     decoded_imm <= $signed({mem_rdata_q[31], mem_rdata_q[7], mem_rdata_q[30:25], mem_rdata_q[11:8], 1'b0});
	   is_sb_sh_sw:
	     decoded_imm <= $signed({mem_rdata_q[31:25], mem_rdata_q[11:7]});
	   default:
	     decoded_imm <= 1'bx;
	 endcase
      end
   end


   // Main State Machine

   localparam cpu_state_trap   = 8'b10000000;
   localparam cpu_state_fetch  = 8'b01000000;
   localparam cpu_state_ld_rs1 = 8'b00100000;
   localparam cpu_state_ld_rs2 = 8'b00010000;
   localparam cpu_state_exec   = 8'b00001000;
   localparam cpu_state_shift  = 8'b00000100;
   localparam cpu_state_stmem  = 8'b00000010;
   localparam cpu_state_ldmem  = 8'b00000001;

   reg [7:0] cpu_state;
   reg [1:0] irq_state;

   `FORMAL_KEEP reg [127:0] ascii_state;

   always @* begin
      ascii_state = "";
      if (cpu_state == cpu_state_trap)   ascii_state = "trap";
      if (cpu_state == cpu_state_fetch)  ascii_state = "fetch";
      if (cpu_state == cpu_state_ld_rs1) ascii_state = "ld_rs1";
      if (cpu_state == cpu_state_ld_rs2) ascii_state = "ld_rs2";
      if (cpu_state == cpu_state_exec)   ascii_state = "exec";
      if (cpu_state == cpu_state_shift)  ascii_state = "shift";
      if (cpu_state == cpu_state_stmem)  ascii_state = "stmem";
      if (cpu_state == cpu_state_ldmem)  ascii_state = "ldmem";
   end

   reg set_mem_do_rinst;
   reg set_mem_do_rdata;
   reg set_mem_do_wdata;

   reg latched_store;
   reg latched_stalu;
   reg latched_branch;
   reg latched_is_lu;
   reg latched_is_lh;
   reg latched_is_lb;
   reg [regindex_bits-1:0] latched_rd;

   reg [31:0]              current_pc;
   assign next_pc = latched_store && latched_branch ? reg_out : reg_next_pc;

   reg [3:0]               pcpi_timeout_counter;
   reg                     pcpi_timeout;

   reg [31:0]              next_irq_pending;
   reg                     do_waitirq;

   reg [31:0]              alu_out, alu_out_q;
   reg                     alu_out_0, alu_out_0_q;
   reg                     alu_wait, alu_wait_2;

   reg [31:0]              alu_add_sub;
   reg                     alu_eq, alu_ltu, alu_lts;

   generate if (TWO_CYCLE_ALU) begin
      always @(posedge clk) begin
	 alu_add_sub <= instr_sub ? reg_op1 - reg_op2 : reg_op1 + reg_op2;
	 alu_eq <= reg_op1 == reg_op2;
	 alu_lts <= $signed(reg_op1) < $signed(reg_op2);
	 alu_ltu <= reg_op1 < reg_op2;
      end
   end else begin
      always @* begin
	 alu_add_sub = instr_sub ? reg_op1 - reg_op2 : reg_op1 + reg_op2;
	 alu_eq = reg_op1 == reg_op2;
	 alu_lts = $signed(reg_op1) < $signed(reg_op2);
	 alu_ltu = reg_op1 < reg_op2;
      end
   end endgenerate

   always @* begin
      alu_out_0 = 'bx;
      (* parallel_case, full_case *)
      case (1'b1)
	instr_beq:
	  alu_out_0 = alu_eq;
	instr_bne:
	  alu_out_0 = !alu_eq;
	instr_bge:
	  alu_out_0 = !alu_lts;
	instr_bgeu:
	  alu_out_0 = !alu_ltu;
	is_slti_blt_slt:
	  alu_out_0 = alu_lts;
	is_sltiu_bltu_sltu:
	  alu_out_0 = alu_ltu;
      endcase

      alu_out = 'bx;
      (* parallel_case, full_case *)
      case (1'b1)
	is_lui_auipc_jal_jalr_addi_add_sub:
	  alu_out = alu_add_sub;
	is_compare:
	  alu_out = alu_out_0;
	instr_xori || instr_xor:
	  alu_out = reg_op1 ^ reg_op2;
	instr_ori || instr_or:
	  alu_out = reg_op1 | reg_op2;
	instr_andi || instr_and:
	  alu_out = reg_op1 & reg_op2;
      endcase
   end

   always @(posedge clk) begin
      trap <= 0;
      reg_sh <= 'bx;
      reg_out <= 'bx;
      set_mem_do_rinst = 0;
      set_mem_do_rdata = 0;
      set_mem_do_wdata = 0;

      alu_out_0_q <= alu_out_0;
      alu_out_q <= alu_out;

      alu_wait <= 0;
      alu_wait_2 <= 0;

      if (WITH_PCPI && CATCH_ILLINSN) begin
	 if (resetn && pcpi_valid && !pcpi_int_wait) begin
	    if (pcpi_timeout_counter)
	      pcpi_timeout_counter <= pcpi_timeout_counter - 1;
	 end else
	   pcpi_timeout_counter <= ~0;
	 pcpi_timeout <= !pcpi_timeout_counter;
      end

      if (ENABLE_COUNTERS)
	count_cycle <= resetn ? count_cycle + 1 : 0;

      next_irq_pending = ENABLE_IRQ ? irq_pending & LATCHED_IRQ : 'bx;

      if (ENABLE_IRQ && ENABLE_IRQ_TIMER && timer) begin
	 if (timer - 1 == 0)
	   next_irq_pending[irq_timer] = 1;
	 timer <= timer - 1;
      end

      if (ENABLE_IRQ) begin
	 next_irq_pending = next_irq_pending | irq;
      end

      decoder_trigger_q <= decoder_trigger;
      decoder_trigger <= mem_do_rinst && mem_done;
      decoder_pseudo_trigger <= 0;
      do_waitirq <= 0;

      if (!resetn) begin
	 reg_pc <= PROGADDR_RESET;
	 reg_next_pc <= PROGADDR_RESET;
	 if (ENABLE_COUNTERS)
	   count_instr <= 0;
	 latched_store <= 0;
	 latched_stalu <= 0;
	 latched_branch <= 0;
	 latched_is_lu <= 0;
	 latched_is_lh <= 0;
	 latched_is_lb <= 0;
	 pcpi_valid <= 0;
	 irq_active <= 0;
	 irq_mask <= ~0;
	 next_irq_pending = 0;
	 irq_state <= 0;
	 eoi <= 0;
	 timer <= 0;
	 cpu_state <= cpu_state_fetch;
      end else
	(* parallel_case, full_case *)
	case (cpu_state)
	  cpu_state_trap: begin
	     trap <= 1;
	  end

	  cpu_state_fetch: begin
	     mem_do_rinst <= !decoder_trigger && !do_waitirq;
	     mem_wordsize <= 0;

	     current_pc = reg_next_pc;

	     (* parallel_case *)
	     case (1'b1)
	       latched_branch: begin
		  current_pc = latched_store ? (latched_stalu ? alu_out_q : reg_out) : reg_next_pc;
		  `debug($display("ST_RD:  %2d 0x%08x, BRANCH 0x%08x", latched_rd, reg_pc + 4, current_pc);)
		  cpuregs[latched_rd] <= reg_pc + 4;
	       end
	       latched_store && !latched_branch: begin
		  `debug($display("ST_RD:  %2d 0x%08x", latched_rd, latched_stalu ? alu_out_q : reg_out);)
		  cpuregs[latched_rd] <= latched_stalu ? alu_out_q : reg_out;
	       end
	       ENABLE_IRQ && irq_state[0]: begin
		  cpuregs[latched_rd] <= current_pc;
		  current_pc = PROGADDR_IRQ;
		  irq_active <= 1;
		  mem_do_rinst <= 1;
	       end
	       ENABLE_IRQ && irq_state[1]: begin
		  eoi <= irq_pending & ~irq_mask;
		  cpuregs[latched_rd] <= irq_pending & ~irq_mask;
		  next_irq_pending = next_irq_pending & irq_mask;
	       end
	     endcase

	     reg_pc <= current_pc;
	     reg_next_pc <= current_pc;

	     latched_store <= 0;
	     latched_stalu <= 0;
	     latched_branch <= 0;
	     latched_is_lu <= 0;
	     latched_is_lh <= 0;
	     latched_is_lb <= 0;
	     latched_rd <= decoded_rd;

	     if (ENABLE_IRQ && ((decoder_trigger && !irq_active && |(irq_pending & ~irq_mask)) || irq_state)) begin
		irq_state <=
			    irq_state == 2'b00 ? 2'b01 :
			    irq_state == 2'b01 ? 2'b10 : 2'b00;
		if (ENABLE_IRQ_QREGS)
		  latched_rd <= irqregs_offset | irq_state[0];
		else
		  latched_rd <= irq_state[0] ? 4 : 3;
	     end else
	       if (ENABLE_IRQ && (decoder_trigger || do_waitirq) && instr_waitirq) begin
		  if (irq_pending) begin
		     latched_store <= 1;
		     reg_out <= irq_pending;
		     reg_next_pc <= current_pc + 4;
		     mem_do_rinst <= 1;
		  end else
		    do_waitirq <= 1;
	       end else
		 if (decoder_trigger) begin
		    `debug($display("-- %-0t", $time);)
		    reg_next_pc <= current_pc + 4;
		    if (ENABLE_COUNTERS)
		      count_instr <= count_instr + 1;
		    if (instr_jal) begin
		       `debug($display("DECODE: 0x%08x jal", current_pc);)
		       mem_do_rinst <= 1;
		       reg_next_pc <= current_pc + decoded_imm_uj;
		       latched_branch <= 1;
		    end else begin
		       mem_do_rinst <= 0;
		       mem_do_prefetch <= !instr_jalr && !instr_retirq;
		       cpu_state <= cpu_state_ld_rs1;
		    end
		 end
	  end

	  cpu_state_ld_rs1: begin
	     reg_op1 <= 'bx;
	     reg_op2 <= 'bx;
	     `debug($display("DECODE: 0x%08x %-0s", reg_pc, ascii_instr ? ascii_instr : "UNKNOWN");)

	     (* parallel_case *)
	     case (1'b1)
	       (CATCH_ILLINSN || WITH_PCPI) && instr_trap: begin
		  if (WITH_PCPI) begin
		     `debug($display("LD_RS1: %2d 0x%08x", decoded_rs1, decoded_rs1 ? cpuregs[decoded_rs1] : 0);)
		     reg_op1 <= decoded_rs1 ? cpuregs[decoded_rs1] : 0;
		     if (ENABLE_REGS_DUALPORT) begin
			pcpi_valid <= 1;
			`debug($display("LD_RS2: %2d 0x%08x", decoded_rs2, decoded_rs2 ? cpuregs[decoded_rs2] : 0);)
			reg_sh <= decoded_rs2 ? cpuregs[decoded_rs2] : 0;
			reg_op2 <= decoded_rs2 ? cpuregs[decoded_rs2] : 0;
			if (pcpi_int_ready) begin
			   mem_do_rinst <= 1;
			   pcpi_valid <= 0;
			   reg_out <= pcpi_int_rd;
			   latched_store <= pcpi_int_wr;
			   cpu_state <= cpu_state_fetch;
			end else
			  if (CATCH_ILLINSN && pcpi_timeout) begin
			     `debug($display("SBREAK OR UNSUPPORTED INSN AT 0x%08x", reg_pc);)
			     if (ENABLE_IRQ && !irq_mask[irq_sbreak] && !irq_active) begin
				next_irq_pending[irq_sbreak] = 1;
				cpu_state <= cpu_state_fetch;
			     end else
			       cpu_state <= cpu_state_trap;
			  end
		     end else begin
			cpu_state <= cpu_state_ld_rs2;
		     end
		  end else begin
		     `debug($display("SBREAK OR UNSUPPORTED INSN AT 0x%08x", reg_pc);)
		     if (ENABLE_IRQ && !irq_mask[irq_sbreak] && !irq_active) begin
			next_irq_pending[irq_sbreak] = 1;
			cpu_state <= cpu_state_fetch;
		     end else
		       cpu_state <= cpu_state_trap;
		  end
	       end
	       ENABLE_COUNTERS && is_rdcycle_rdcycleh_rdinstr_rdinstrh: begin
		  (* parallel_case, full_case *)
		  case (1'b1)
		    instr_rdcycle:
		      reg_out <= count_cycle[31:0];
		    instr_rdcycleh:
		      reg_out <= count_cycle[63:32];
		    instr_rdinstr:
		      reg_out <= count_instr[31:0];
		    instr_rdinstrh:
		      reg_out <= count_instr[63:32];
		  endcase
		  latched_store <= 1;
		  cpu_state <= cpu_state_fetch;
	       end
	       is_lui_auipc_jal: begin
		  reg_op1 <= instr_lui ? 0 : reg_pc;
		  reg_op2 <= decoded_imm;
		  if (TWO_CYCLE_ALU)
		    alu_wait <= 1;
		  else
		    mem_do_rinst <= mem_do_prefetch;
		  cpu_state <= cpu_state_exec;
	       end
	       ENABLE_IRQ && ENABLE_IRQ_QREGS && instr_getq: begin
		  `debug($display("LD_RS1: %2d 0x%08x", decoded_rs1, decoded_rs1 ? cpuregs[decoded_rs1] : 0);)
		  reg_out <= decoded_rs1 ? cpuregs[decoded_rs1] : 0;
		  latched_store <= 1;
		  cpu_state <= cpu_state_fetch;
	       end
	       ENABLE_IRQ && ENABLE_IRQ_QREGS && instr_setq: begin
		  `debug($display("LD_RS1: %2d 0x%08x", decoded_rs1, decoded_rs1 ? cpuregs[decoded_rs1] : 0);)
		  reg_out <= decoded_rs1 ? cpuregs[decoded_rs1] : 0;
		  latched_rd <= latched_rd | irqregs_offset;
		  latched_store <= 1;
		  cpu_state <= cpu_state_fetch;
	       end
	       ENABLE_IRQ && instr_retirq: begin
		  eoi <= 0;
		  irq_active <= 0;
		  latched_branch <= 1;
		  latched_store <= 1;
		  `debug($display("LD_RS1: %2d 0x%08x", decoded_rs1, decoded_rs1 ? cpuregs[decoded_rs1] : 0);)
		  reg_out <= decoded_rs1 ? cpuregs[decoded_rs1] : 0;
		  cpu_state <= cpu_state_fetch;
	       end
	       ENABLE_IRQ && instr_maskirq: begin
		  latched_store <= 1;
		  reg_out <= irq_mask;
		  `debug($display("LD_RS1: %2d 0x%08x", decoded_rs1, decoded_rs1 ? cpuregs[decoded_rs1] : 0);)
		  irq_mask <= (decoded_rs1 ? cpuregs[decoded_rs1] : 0) | MASKED_IRQ;
		  cpu_state <= cpu_state_fetch;
	       end
	       ENABLE_IRQ && ENABLE_IRQ_TIMER && instr_timer: begin
		  latched_store <= 1;
		  reg_out <= timer;
		  `debug($display("LD_RS1: %2d 0x%08x", decoded_rs1, decoded_rs1 ? cpuregs[decoded_rs1] : 0);)
		  timer <= decoded_rs1 ? cpuregs[decoded_rs1] : 0;
		  cpu_state <= cpu_state_fetch;
	       end
	       is_lb_lh_lw_lbu_lhu: begin
		  `debug($display("LD_RS1: %2d 0x%08x", decoded_rs1, decoded_rs1 ? cpuregs[decoded_rs1] : 0);)
		  reg_op1 <= decoded_rs1 ? cpuregs[decoded_rs1] : 0;
		  cpu_state <= cpu_state_ldmem;
		  mem_do_rinst <= 1;
	       end
	       is_slli_srli_srai: begin
		  `debug($display("LD_RS1: %2d 0x%08x", decoded_rs1, decoded_rs1 ? cpuregs[decoded_rs1] : 0);)
		  reg_op1 <= decoded_rs1 ? cpuregs[decoded_rs1] : 0;
		  reg_sh <= decoded_rs2;
		  cpu_state <= cpu_state_shift;
	       end
	       is_jalr_addi_slti_sltiu_xori_ori_andi: begin
		  `debug($display("LD_RS1: %2d 0x%08x", decoded_rs1, decoded_rs1 ? cpuregs[decoded_rs1] : 0);)
		  reg_op1 <= decoded_rs1 ? cpuregs[decoded_rs1] : 0;
		  reg_op2 <= decoded_imm;
		  if (TWO_CYCLE_ALU)
		    alu_wait <= 1;
		  else
		    mem_do_rinst <= mem_do_prefetch;
		  cpu_state <= cpu_state_exec;
	       end
	       default: begin
		  `debug($display("LD_RS1: %2d 0x%08x", decoded_rs1, decoded_rs1 ? cpuregs[decoded_rs1] : 0);)
		  reg_op1 <= decoded_rs1 ? cpuregs[decoded_rs1] : 0;
		  if (ENABLE_REGS_DUALPORT) begin
		     `debug($display("LD_RS2: %2d 0x%08x", decoded_rs2, decoded_rs2 ? cpuregs[decoded_rs2] : 0);)
		     reg_sh <= decoded_rs2 ? cpuregs[decoded_rs2] : 0;
		     reg_op2 <= decoded_rs2 ? cpuregs[decoded_rs2] : 0;
		     (* parallel_case *)
		     case (1'b1)
		       is_sb_sh_sw: begin
			  cpu_state <= cpu_state_stmem;
			  mem_do_rinst <= 1;
		       end
		       is_sll_srl_sra: begin
			  cpu_state <= cpu_state_shift;
		       end
		       default: begin
			  if (TWO_CYCLE_ALU || (TWO_CYCLE_COMPARE && is_beq_bne_blt_bge_bltu_bgeu)) begin
			     alu_wait_2 <= TWO_CYCLE_ALU && (TWO_CYCLE_COMPARE && is_beq_bne_blt_bge_bltu_bgeu);
			     alu_wait <= 1;
			  end else
			    mem_do_rinst <= mem_do_prefetch;
			  cpu_state <= cpu_state_exec;
		       end
		     endcase
		  end else
		    cpu_state <= cpu_state_ld_rs2;
	       end
	     endcase
	  end

	  cpu_state_ld_rs2: begin
	     `debug($display("LD_RS2: %2d 0x%08x", decoded_rs2, decoded_rs2 ? cpuregs[decoded_rs2] : 0);)
	     reg_sh <= decoded_rs2 ? cpuregs[decoded_rs2] : 0;
	     reg_op2 <= decoded_rs2 ? cpuregs[decoded_rs2] : 0;

	     (* parallel_case *)
	     case (1'b1)
	       WITH_PCPI && instr_trap: begin
		  pcpi_valid <= 1;
		  if (pcpi_int_ready) begin
		     mem_do_rinst <= 1;
		     pcpi_valid <= 0;
		     reg_out <= pcpi_int_rd;
		     latched_store <= pcpi_int_wr;
		     cpu_state <= cpu_state_fetch;
		  end else
		    if (CATCH_ILLINSN && pcpi_timeout) begin
		       `debug($display("SBREAK OR UNSUPPORTED INSN AT 0x%08x", reg_pc);)
		       if (ENABLE_IRQ && !irq_mask[irq_sbreak] && !irq_active) begin
			  next_irq_pending[irq_sbreak] = 1;
			  cpu_state <= cpu_state_fetch;
		       end else
			 cpu_state <= cpu_state_trap;
		    end
	       end
	       is_sb_sh_sw: begin
		  cpu_state <= cpu_state_stmem;
		  mem_do_rinst <= 1;
	       end
	       is_sll_srl_sra: begin
		  cpu_state <= cpu_state_shift;
	       end
	       default: begin
		  if (TWO_CYCLE_ALU || (TWO_CYCLE_COMPARE && is_beq_bne_blt_bge_bltu_bgeu)) begin
		     alu_wait_2 <= TWO_CYCLE_ALU && (TWO_CYCLE_COMPARE && is_beq_bne_blt_bge_bltu_bgeu);
		     alu_wait <= 1;
		  end else
		    mem_do_rinst <= mem_do_prefetch;
		  cpu_state <= cpu_state_exec;
	       end
	     endcase
	  end

	  cpu_state_exec: begin
	     latched_store <= TWO_CYCLE_COMPARE ? alu_out_0_q : alu_out_0;
	     latched_branch <= TWO_CYCLE_COMPARE ? alu_out_0_q : alu_out_0;
	     reg_out <= reg_pc + decoded_imm;
	     if ((TWO_CYCLE_ALU || TWO_CYCLE_COMPARE) && (alu_wait || alu_wait_2)) begin
		mem_do_rinst <= mem_do_prefetch && !alu_wait_2;
		alu_wait <= alu_wait_2;
	     end else
	       if (is_beq_bne_blt_bge_bltu_bgeu) begin
		  latched_rd <= 0;
		  if (mem_done)
		    cpu_state <= cpu_state_fetch;
		  if (TWO_CYCLE_COMPARE ? alu_out_0_q : alu_out_0) begin
		     decoder_trigger <= 0;
		     set_mem_do_rinst = 1;
		  end
	       end else begin
		  latched_branch <= instr_jalr;
		  latched_store <= 1;
		  latched_stalu <= 1;
		  cpu_state <= cpu_state_fetch;
	       end
	  end

	  cpu_state_shift: begin
	     latched_store <= 1;
	     if (reg_sh == 0) begin
		reg_out <= reg_op1;
		mem_do_rinst <= mem_do_prefetch;
		cpu_state <= cpu_state_fetch;
	     end else if (TWO_STAGE_SHIFT && reg_sh >= 4) begin
		(* parallel_case, full_case *)
		case (1'b1)
		  instr_slli || instr_sll: reg_op1 <= reg_op1 << 4;
		  instr_srli || instr_srl: reg_op1 <= reg_op1 >> 4;
		  instr_srai || instr_sra: reg_op1 <= $signed(reg_op1) >>> 4;
		endcase
		reg_sh <= reg_sh - 4;
	     end else begin
		(* parallel_case, full_case *)
		case (1'b1)
		  instr_slli || instr_sll: reg_op1 <= reg_op1 << 1;
		  instr_srli || instr_srl: reg_op1 <= reg_op1 >> 1;
		  instr_srai || instr_sra: reg_op1 <= $signed(reg_op1) >>> 1;
		endcase
		reg_sh <= reg_sh - 1;
	     end
	  end

	  cpu_state_stmem: begin
	     if (!mem_do_prefetch || mem_done) begin
		if (!mem_do_wdata) begin
		   (* parallel_case, full_case *)
		   case (1'b1)
		     instr_sb: mem_wordsize <= 2;
		     instr_sh: mem_wordsize <= 1;
		     instr_sw: mem_wordsize <= 0;
		   endcase
		   reg_op1 <= reg_op1 + decoded_imm;
		   set_mem_do_wdata = 1;
		end
		if (!mem_do_prefetch && mem_done) begin
		   cpu_state <= cpu_state_fetch;
		   decoder_trigger <= 1;
		   decoder_pseudo_trigger <= 1;
		end
	     end
	  end

	  cpu_state_ldmem: begin
	     latched_store <= 1;
	     if (!mem_do_prefetch || mem_done) begin
		if (!mem_do_rdata) begin
		   (* parallel_case, full_case *)
		   case (1'b1)
		     instr_lb || instr_lbu: mem_wordsize <= 2;
		     instr_lh || instr_lhu: mem_wordsize <= 1;
		     instr_lw: mem_wordsize <= 0;
		   endcase
		   latched_is_lu <= is_lbu_lhu_lw;
		   latched_is_lh <= instr_lh;
		   latched_is_lb <= instr_lb;
		   reg_op1 <= reg_op1 + decoded_imm;
		   set_mem_do_rdata = 1;
		end
		if (!mem_do_prefetch && mem_done) begin
		   (* parallel_case, full_case *)
		   case (1'b1)
		     latched_is_lu: reg_out <= mem_rdata_word;
		     latched_is_lh: reg_out <= $signed(mem_rdata_word[15:0]);
		     latched_is_lb: reg_out <= $signed(mem_rdata_word[7:0]);
		   endcase
		   decoder_trigger <= 1;
		   decoder_pseudo_trigger <= 1;
		   cpu_state <= cpu_state_fetch;
		end
	     end
	  end
	endcase

      if (CATCH_MISALIGN && resetn && (mem_do_rdata || mem_do_wdata)) begin
	 if (mem_wordsize == 0 && reg_op1[1:0] != 0) begin
	    `debug($display("MISALIGNED WORD: 0x%08x", reg_op1);)
	    if (ENABLE_IRQ && !irq_mask[irq_buserror] && !irq_active) begin
	       next_irq_pending[irq_buserror] = 1;
	    end else
	      cpu_state <= cpu_state_trap;
	 end
	 if (mem_wordsize == 1 && reg_op1[0] != 0) begin
	    `debug($display("MISALIGNED HALFWORD: 0x%08x", reg_op1);)
	    if (ENABLE_IRQ && !irq_mask[irq_buserror] && !irq_active) begin
	       next_irq_pending[irq_buserror] = 1;
	    end else
	      cpu_state <= cpu_state_trap;
	 end
      end
      if (CATCH_MISALIGN && resetn && mem_do_rinst && reg_pc[1:0] != 0) begin
	 `debug($display("MISALIGNED INSTRUCTION: 0x%08x", reg_pc);)
	 if (ENABLE_IRQ && !irq_mask[irq_buserror] && !irq_active) begin
	    next_irq_pending[irq_buserror] = 1;
	 end else
	   cpu_state <= cpu_state_trap;
      end

      if (!resetn || mem_done) begin
	 mem_do_prefetch <= 0;
	 mem_do_rinst <= 0;
	 mem_do_rdata <= 0;
	 mem_do_wdata <= 0;
      end

      if (set_mem_do_rinst)
	mem_do_rinst <= 1;
      if (set_mem_do_rdata)
	mem_do_rdata <= 1;
      if (set_mem_do_wdata)
	mem_do_wdata <= 1;

      irq_pending <= next_irq_pending & ~MASKED_IRQ;

      reg_pc[1:0] <= 0;
      reg_next_pc[1:0] <= 0;
      current_pc = 'bx;
   end


   // Formal Verification
`ifdef FORMAL
   reg [3:0] cycle = 0;
   always @(posedge clk)
     if (~&cycle) cycle <= cycle + 1;

   reg [4:0] last_mem_ready;
   always @(posedge clk)
     last_mem_ready <= {last_mem_ready, mem_ready};
   assume property (|last_mem_ready);

   reg       ok;
   always @* begin
      assume (resetn == |cycle);
      if (cycle) begin
	 // instruction fetches are read-only
	 if (mem_valid && mem_instr)
	   assert (mem_wstrb == 0);

	 // cpu_state must be valid
	 ok = 0;
	 if (cpu_state == cpu_state_trap)   ok = 1;
	 if (cpu_state == cpu_state_fetch)  ok = 1;
	 if (cpu_state == cpu_state_ld_rs1) ok = 1;
	 if (cpu_state == cpu_state_ld_rs2) ok = ENABLE_REGS_DUALPORT;
	 if (cpu_state == cpu_state_exec)   ok = 1;
	 if (cpu_state == cpu_state_shift)  ok = 1;
	 if (cpu_state == cpu_state_stmem)  ok = 1;
	 if (cpu_state == cpu_state_ldmem)  ok = 1;
	 assert (ok);
      end
   end
`endif
endmodule


/***************************************************************
 * picorv32_pcpi_mul
 ***************************************************************/

module picorv32_pcpi_mul #(
	                   parameter STEPS_AT_ONCE = 1,
	                   parameter CARRY_CHAIN = 4
                           ) (
	                      input             clk, resetn,

	                      input             pcpi_valid,
	                      input [31:0]      pcpi_insn,
	                      input [31:0]      pcpi_rs1,
	                      input [31:0]      pcpi_rs2,
	                      output reg        pcpi_wr,
	                      output reg [31:0] pcpi_rd,
	                      output reg        pcpi_wait,
	                      output reg        pcpi_ready
                              );
   reg                                          instr_mul, instr_mulh, instr_mulhsu, instr_mulhu;
   wire                                         instr_any_mul = |{instr_mul, instr_mulh, instr_mulhsu, instr_mulhu};
   wire                                         instr_any_mulh = |{instr_mulh, instr_mulhsu, instr_mulhu};
   wire                                         instr_rs1_signed = |{instr_mulh, instr_mulhsu};
   wire                                         instr_rs2_signed = |{instr_mulh};

   reg                                          pcpi_wait_q;
   wire                                         mul_start = pcpi_wait && !pcpi_wait_q;

   always @(posedge clk) begin
      instr_mul <= 0;
      instr_mulh <= 0;
      instr_mulhsu <= 0;
      instr_mulhu <= 0;

      if (resetn && pcpi_valid && pcpi_insn[6:0] == 7'b0110011 && pcpi_insn[31:25] == 7'b0000001) begin
	 case (pcpi_insn[14:12])
	   3'b000: instr_mul <= 1;
	   3'b001: instr_mulh <= 1;
	   3'b010: instr_mulhsu <= 1;
	   3'b011: instr_mulhu <= 1;
	 endcase
      end

      pcpi_wait <= instr_any_mul;
      pcpi_wait_q <= pcpi_wait;
   end

   reg [63:0] rs1, rs2, rd, rdx;
   reg [63:0] next_rs1, next_rs2, this_rs2;
   reg [63:0] next_rd, next_rdx, next_rdt;
   reg [6:0]  mul_counter;
   reg        mul_waiting;
   reg        mul_finish;
   integer    i, j;

   // carry save accumulator
   always @* begin
      next_rd = rd;
      next_rdx = rdx;
      next_rs1 = rs1;
      next_rs2 = rs2;

      for (i = 0; i < STEPS_AT_ONCE; i=i+1) begin
	 this_rs2 = next_rs1[0] ? next_rs2 : 0;
	 if (CARRY_CHAIN == 0) begin
	    next_rdt = next_rd ^ next_rdx ^ this_rs2;
	    next_rdx = ((next_rd & next_rdx) | (next_rd & this_rs2) | (next_rdx & this_rs2)) << 1;
	    next_rd = next_rdt;
	 end else begin
	    next_rdt = 0;
	    for (j = 0; j < 64; j = j + CARRY_CHAIN)
	      {next_rdt[j+CARRY_CHAIN-1], next_rd[j +: CARRY_CHAIN]} =
		     next_rd[j +: CARRY_CHAIN] + next_rdx[j +: CARRY_CHAIN] + this_rs2[j +: CARRY_CHAIN];
	    next_rdx = next_rdt << 1;
	 end
	 next_rs1 = next_rs1 >> 1;
	 next_rs2 = next_rs2 << 1;
      end
   end

   always @(posedge clk) begin
      mul_finish <= 0;
      if (!resetn) begin
	 mul_waiting <= 1;
      end else
	if (mul_waiting) begin
	   if (instr_rs1_signed)
	     rs1 <= $signed(pcpi_rs1);
	   else
	     rs1 <= $unsigned(pcpi_rs1);

	   if (instr_rs2_signed)
	     rs2 <= $signed(pcpi_rs2);
	   else
	     rs2 <= $unsigned(pcpi_rs2);

	   rd <= 0;
	   rdx <= 0;
	   mul_counter <= (instr_any_mulh ? 63 - STEPS_AT_ONCE : 31 - STEPS_AT_ONCE);
	   mul_waiting <= !mul_start;
	end else begin
	   rd <= next_rd;
	   rdx <= next_rdx;
	   rs1 <= next_rs1;
	   rs2 <= next_rs2;

	   mul_counter <= mul_counter - STEPS_AT_ONCE;
	   if (mul_counter[6]) begin
	      mul_finish <= 1;
	      mul_waiting <= 1;
	   end
	end
   end

   always @(posedge clk) begin
      pcpi_wr <= 0;
      pcpi_ready <= 0;
      if (mul_finish) begin
	 pcpi_wr <= 1;
	 pcpi_ready <= 1;
	 pcpi_rd <= instr_any_mulh ? rd >> 32 : rd;
      end
   end
endmodule


/***************************************************************
 * picorv32_axi
 ***************************************************************/

module picorv32_axi #(
	              parameter [ 0:0] ENABLE_COUNTERS = 1,
	              parameter [ 0:0] ENABLE_REGS_16_31 = 1,
	              parameter [ 0:0] ENABLE_REGS_DUALPORT = 1,
	              parameter [ 0:0] TWO_STAGE_SHIFT = 1,
	              parameter [ 0:0] TWO_CYCLE_COMPARE = 0,
	              parameter [ 0:0] TWO_CYCLE_ALU = 0,
	              parameter [ 0:0] CATCH_MISALIGN = 1,
	              parameter [ 0:0] CATCH_ILLINSN = 1,
	              parameter [ 0:0] ENABLE_PCPI = 0,
	              parameter [ 0:0] ENABLE_MUL = 0,
	              parameter [ 0:0] ENABLE_IRQ = 0,
	              parameter [ 0:0] ENABLE_IRQ_QREGS = 1,
	              parameter [ 0:0] ENABLE_IRQ_TIMER = 1,
	              parameter [31:0] MASKED_IRQ = 32'h 0000_0000,
	              parameter [31:0] LATCHED_IRQ = 32'h ffff_ffff,
	              parameter [31:0] PROGADDR_RESET = 32'h 0000_0000,
	              parameter [31:0] PROGADDR_IRQ = 32'h 0000_0010
                      ) (
	                 input         clk, resetn,
	                 output        trap,

	                 // AXI4-lite master memory interface

	                 output        mem_axi_awvalid,
	                 input         mem_axi_awready,
	                 output [31:0] mem_axi_awaddr,
	                 output [ 2:0] mem_axi_awprot,

	                 output        mem_axi_wvalid,
	                 input         mem_axi_wready,
	                 output [31:0] mem_axi_wdata,
	                 output [ 3:0] mem_axi_wstrb,

	                 input         mem_axi_bvalid,
	                 output        mem_axi_bready,

	                 output        mem_axi_arvalid,
	                 input         mem_axi_arready,
	                 output [31:0] mem_axi_araddr,
	                 output [ 2:0] mem_axi_arprot,

	                 input         mem_axi_rvalid,
	                 output        mem_axi_rready,
	                 input [31:0]  mem_axi_rdata,

	                 // Pico Co-Processor Interface (PCPI)
	                 output        pcpi_valid,
	                 output [31:0] pcpi_insn,
	                 output [31:0] pcpi_rs1,
	                 output [31:0] pcpi_rs2,
	                 input         pcpi_wr,
	                 input [31:0]  pcpi_rd,
	                 input         pcpi_wait,
	                 input         pcpi_ready,

	                 // IRQ interface
	                 input [31:0]  irq,
	                 output [31:0] eoi
                         );
   wire                                mem_valid;
   wire [31:0]                         mem_addr;
   wire [31:0]                         mem_wdata;
   wire [ 3:0]                         mem_wstrb;
   wire                                mem_instr;
   wire                                mem_ready;
   wire [31:0]                         mem_rdata;

   picorv32_axi_adapter axi_adapter (
		                     .clk            (clk            ),
		                     .resetn         (resetn         ),
		                     .mem_axi_awvalid(mem_axi_awvalid),
		                     .mem_axi_awready(mem_axi_awready),
		                     .mem_axi_awaddr (mem_axi_awaddr ),
		                     .mem_axi_awprot (mem_axi_awprot ),
		                     .mem_axi_wvalid (mem_axi_wvalid ),
		                     .mem_axi_wready (mem_axi_wready ),
		                     .mem_axi_wdata  (mem_axi_wdata  ),
		                     .mem_axi_wstrb  (mem_axi_wstrb  ),
		                     .mem_axi_bvalid (mem_axi_bvalid ),
		                     .mem_axi_bready (mem_axi_bready ),
		                     .mem_axi_arvalid(mem_axi_arvalid),
		                     .mem_axi_arready(mem_axi_arready),
		                     .mem_axi_araddr (mem_axi_araddr ),
		                     .mem_axi_arprot (mem_axi_arprot ),
		                     .mem_axi_rvalid (mem_axi_rvalid ),
		                     .mem_axi_rready (mem_axi_rready ),
		                     .mem_axi_rdata  (mem_axi_rdata  ),
		                     .mem_valid      (mem_valid      ),
		                     .mem_instr      (mem_instr      ),
		                     .mem_ready      (mem_ready      ),
		                     .mem_addr       (mem_addr       ),
		                     .mem_wdata      (mem_wdata      ),
		                     .mem_wstrb      (mem_wstrb      ),
		                     .mem_rdata      (mem_rdata      )
	                             );

   picorv32 #(
	      .ENABLE_COUNTERS     (ENABLE_COUNTERS     ),
	      .ENABLE_REGS_16_31   (ENABLE_REGS_16_31   ),
	      .ENABLE_REGS_DUALPORT(ENABLE_REGS_DUALPORT),
	      .TWO_STAGE_SHIFT     (TWO_STAGE_SHIFT     ),
	      .TWO_CYCLE_COMPARE   (TWO_CYCLE_COMPARE   ),
	      .TWO_CYCLE_ALU       (TWO_CYCLE_ALU       ),
	      .CATCH_MISALIGN      (CATCH_MISALIGN      ),
	      .CATCH_ILLINSN       (CATCH_ILLINSN       ),
	      .ENABLE_PCPI         (ENABLE_PCPI         ),
	      .ENABLE_MUL          (ENABLE_MUL          ),
	      .ENABLE_IRQ          (ENABLE_IRQ          ),
	      .ENABLE_IRQ_QREGS    (ENABLE_IRQ_QREGS    ),
	      .ENABLE_IRQ_TIMER    (ENABLE_IRQ_TIMER    ),
	      .MASKED_IRQ          (MASKED_IRQ          ),
	      .LATCHED_IRQ         (LATCHED_IRQ         ),
	      .PROGADDR_RESET      (PROGADDR_RESET      ),
	      .PROGADDR_IRQ        (PROGADDR_IRQ        )
	      ) picorv32_core (
		               .clk      (clk   ),
		               .resetn   (resetn),
		               .trap     (trap  ),

		               .mem_valid(mem_valid),
		               .mem_addr (mem_addr ),
		               .mem_wdata(mem_wdata),
		               .mem_wstrb(mem_wstrb),
		               .mem_instr(mem_instr),
		               .mem_ready(mem_ready),
		               .mem_rdata(mem_rdata),

		               .pcpi_valid(pcpi_valid),
		               .pcpi_insn (pcpi_insn ),
		               .pcpi_rs1  (pcpi_rs1  ),
		               .pcpi_rs2  (pcpi_rs2  ),
		               .pcpi_wr   (pcpi_wr   ),
		               .pcpi_rd   (pcpi_rd   ),
		               .pcpi_wait (pcpi_wait ),
		               .pcpi_ready(pcpi_ready),

		               .irq(irq),
		               .eoi(eoi)
	                       );
endmodule


/***************************************************************
 * picorv32_axi_adapter
 ***************************************************************/

module picorv32_axi_adapter (
	                     input         clk, resetn,

	                     // AXI4-lite master memory interface

	                     output        mem_axi_awvalid,
	                     input         mem_axi_awready,
	                     output [31:0] mem_axi_awaddr,
	                     output [ 2:0] mem_axi_awprot,

	                     output        mem_axi_wvalid,
	                     input         mem_axi_wready,
	                     output [31:0] mem_axi_wdata,
	                     output [ 3:0] mem_axi_wstrb,

	                     input         mem_axi_bvalid,
	                     output        mem_axi_bready,

	                     output        mem_axi_arvalid,
	                     input         mem_axi_arready,
	                     output [31:0] mem_axi_araddr,
	                     output [ 2:0] mem_axi_arprot,

	                     input         mem_axi_rvalid,
	                     output        mem_axi_rready,
	                     input [31:0]  mem_axi_rdata,

	                     // Native PicoRV32 memory interface

	                     input         mem_valid,
	                     input         mem_instr,
	                     output        mem_ready,
	                     input [31:0]  mem_addr,
	                     input [31:0]  mem_wdata,
	                     input [ 3:0]  mem_wstrb,
	                     output [31:0] mem_rdata
                             );
   reg                                     ack_awvalid;
   reg                                     ack_arvalid;
   reg                                     ack_wvalid;

   assign mem_axi_awvalid = mem_valid && |mem_wstrb && !ack_awvalid;
   assign mem_axi_awaddr = mem_addr;
   assign mem_axi_awprot = 0;

   assign mem_axi_arvalid = mem_valid && !mem_wstrb && !ack_arvalid;
   assign mem_axi_araddr = mem_addr;
   assign mem_axi_arprot = mem_instr ? 3'b100 : 3'b000;

   assign mem_axi_wvalid = mem_valid && |mem_wstrb && !ack_wvalid;
   assign mem_axi_wdata = mem_wdata;
   assign mem_axi_wstrb = mem_wstrb;

   assign mem_ready = mem_axi_bvalid || mem_axi_rvalid;
   assign mem_axi_bready = mem_valid && |mem_wstrb;
   assign mem_axi_rready = mem_valid && !mem_wstrb;
   assign mem_rdata = mem_axi_rdata;

   always @(posedge clk) begin
      if (!resetn) begin
	 ack_awvalid <= 0;
      end else begin
	 if (mem_axi_awready && mem_axi_awvalid)
	   ack_awvalid <= 1;
	 if (mem_axi_arready && mem_axi_arvalid)
	   ack_arvalid <= 1;
	 if (mem_axi_wready && mem_axi_wvalid)
	   ack_wvalid <= 1;
	 if (!mem_valid) begin
	    ack_awvalid <= 0;
	    ack_arvalid <= 0;
	    ack_wvalid <= 0;
	 end
      end
   end
endmodule
